
module J_K_FF(
input J,K,clk,
output reg Q,
output Qbar);
always@(posedge clk)
begin 
case ({J,K})
2'b00 : Q <= Q;
2'b01 : Q <= 1'b0;
2'b10 : Q <= 1'b1;
2'b11 : Q <= ~Q;
endcase
end
assign Qbar = ~Q;
endmodule
